** Profile: "SCHEMATIC1-Simulare"  [ f:\facultate\an2\semestrul 2\tehnici cad\proiect\proiect-pspicefiles\schematic1\simulare.sim ] 

** Creating circuit file "Simulare.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../led_violet.lib" 
.LIB "../../../led_verde.lib" 
.LIB "../../../led_rosu.lib" 
.LIB "../../../led_galben.lib" 
.LIB "../../../led_albastru.lib" 
.LIB "../../../led_alb.lib" 
* From [PSPICE NETLIST] section of C:\Users\Mihai\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 0.1m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
